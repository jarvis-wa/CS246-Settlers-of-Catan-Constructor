2
51 57 52 47 43 r h 47 B 53 B
0 1 0 1 2 r h 42 B 45 B
5 6 5 5 4 r h 30 B 33 B
10 10 10 10 20 r h 8 B 26 B
0 3 1 10 3 5 1 4 5 7 3 10 2 11 0 3 3 8 0 2 0 6 1 8 4 12 1 5 4 11 2 4 4 6 2 9 2 9
4
